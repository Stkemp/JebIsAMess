`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/24/2018 02:54:05 AM
// Design Name: 
// Module Name: multiplier_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module multiplier_tb(

    );
    reg [3:0] m,q;
    wire [7:0] p;
    
    multiplier UUT( .m(m), .p(p), .q(q)); 
    
    initial
    begin
    m=0;
    q=0;
    #20;
    q[0]=0; // q is 1
    m[0]=1; // m is 1
    #20;
    m[0]=0;
    m[1]=1; //2
    #20;
    m[0]=1; //3
    #20;
    m[0]=0; m[1]=0; m[2]=1; //4
    #20;
    m[0]=1; //5
    #20;
    m[0]=0; m[1]=1; //6
    #20;
    m[0]=1; //7 
    #20;
    m[0]=0; m[1]=0; m[2]=0; m[3]=1; //8
    #20;
    m[0]=1; //9
    #20;
    m[0]=0; m[1]=1; //10
    #20;
    m[0]=1; //11
    #20;
    m[0]=0; m[1]=0; m[2]=1; //12
    #20;
    m[0]=1; //13
    #20;
    m[0]=0; m[1]=1; //14
    #20;
    m[0]=1; //15
    #20; //now testing q
    m=0; 
     q[0]=1; // q is 1
       #20;
       q[0]=0;
       q[1]=1; //2
       #20;
       q[0]=1; //3
       #20;
       q[0]=0; q[1]=0; q[2]=1; //4
       #20;
       q[0]=1; //5
       #20;
       q[0]=0; q[1]=1; //6
       #20;
       q[0]=1; //7 
       #20;
       q[0]=0; q[1]=0; q[2]=0; q[3]=1; //8
       #20;
       q[0]=1; //9
       #20;
       q[0]=0; q[1]=1; //10
       #20;
       q[0]=1; //11
       #20;
       q[0]=0; q[1]=0; q[2]=1; //12
       #20;
       q[0]=1; //13
       #20;
       q[0]=0; q[1]=1; //14
       #20;
       q[0]=1; //15
       #20; //now testing squares
       q=0;
       #20; 
       q[0]=1; // q is 1
        m[0]=1; // m is 1
             #20;
             q[0]=0;
             q[1]=1; //2
              m[0]=0;
                m[1]=1; //2
             #20;
             q[0]=1; //3
             m[0]=1; //3
             #20;
             q[0]=0; q[1]=0; q[2]=1; //4
             m[0]=0; m[1]=0; m[2]=1; //4
             #20;
             q[0]=1; //5
             m[0]=1; //5
             #20;
             q[0]=0; q[1]=1; //6
               m[0]=0; m[1]=1; //6
             #20;
             q[0]=1; //7 
              m[0]=1; //7
             #20;
             q[0]=0; q[1]=0; q[2]=0; q[3]=1; //8
             m[0]=0; m[1]=0; m[2]=0; m[3]=1; //8
             #20;
             q[0]=1; //9
              m[0]=1; //9
             #20;
             q[0]=0; q[1]=1; //10
             m[0]=0; m[1]=1; //10
             #20;
             q[0]=1; //11
             m[0]=1;
             #20;
             q[0]=0; q[1]=0; q[2]=1; //12
              m[0]=0; m[1]=0; m[2]=1;
             #20;
             q[0]=1; //13
             m[0]=1;
             #20;
             q[0]=0; q[1]=1; //14
              m[0]=0; m[1]=1; //14
             #20;
             q[0]=1; //15
              m[0]=1;
       
         
    end
endmodule
